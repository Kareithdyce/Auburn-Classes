    Mac OS X            	   2   �      �                                      ATTR       �   �   <                  �   <  com.apple.quarantine q/0081;5c4cc1f8;Chrome;3FE13A29-2365-431D-8AB6-A5803015316F 