    Mac OS X            	   2   �      �                                      ATTR       �   �   <                  �   <  com.apple.quarantine q/0081;5c6f180b;Chrome;742A8ABD-7BAF-47D5-B370-0E9944A5CE61 