    Mac OS X            	   2   �      �                                      ATTR       �   �   <                  �   <  com.apple.quarantine q/0081;5ca655e5;Chrome;5B9A1291-17DD-4F27-AD4B-0EE99F4CDDD5 